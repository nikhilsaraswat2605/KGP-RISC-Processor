`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// name - Amit Kumar, Nikhil Saraswat
// Roll- 20CS30003, 20CS10039
// COA - KGP_RISC
//////////////////////////////////////////////////////////////////////////////////
module Diff(rs, rt, out
    );
	 input [31:0] rs;
	 input [31:0] rt;
	 output reg [31:0] out;
	 reg [31:0] temp;
	 always @(*) begin
		temp = rs ^ rt;
		temp = temp ^ (temp-1);
	 
		case(temp)
			32'b1 : out = 32'd1;
			32'b11 : out = 32'd2;
			32'b111 : out = 32'd3;
			32'b1111 : out = 32'd4;
			
			32'b11111 : out = 32'd5;
			32'b111111 : out = 32'd6;
			32'b1111111 : out = 32'd7;
			32'b11111111 : out = 32'd8;
			
			32'b111111111 : out = 32'd9;
			32'b1111111111 : out = 32'd10;
			32'b11111111111 : out = 32'd11;
			32'b111111111111 : out = 32'd12;
			
			32'b1111111111111 : out = 32'd13;
			32'b11111111111111 : out = 32'd14;
			32'b111111111111111 : out = 32'd15;
			32'b1111111111111111 : out = 32'd16;
			
			
			32'b11111111111111111 : out = 32'd17;
			32'b111111111111111111 : out = 32'd18;
			32'b1111111111111111111 : out = 32'd19;
			32'b11111111111111111111 : out = 32'd20;
			
			32'b111111111111111111111 : out = 32'd21;
			32'b1111111111111111111111 : out = 32'd22;
			32'b11111111111111111111111 : out = 32'd23;
			32'b111111111111111111111111 : out = 32'd24;
			
			32'b1111111111111111111111111 : out = 32'd25;
			32'b11111111111111111111111111 : out = 32'd26;
			32'b111111111111111111111111111 : out = 32'd27;
			32'b1111111111111111111111111111 : out = 32'd28;
			
			32'b11111111111111111111111111111 : out = 32'd29;
			32'b111111111111111111111111111111 : out = 32'd30;
			32'b1111111111111111111111111111111 : out = 32'd31;
			32'b11111111111111111111111111111111 : out = 32'd32;

			default : out = 32'd33;
		endcase
	 end

endmodule
